LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY sl2 IS -- shift left by 2
    PORT (
        a : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        y : OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END;
ARCHITECTURE behave OF sl2 IS
BEGIN
    y <= a(29 DOWNTO 0) & "00";
END;